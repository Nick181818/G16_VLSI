module top_module( 
    input a,b,c,
    output reg w,x,y,z );
    assign w=a;
    assign x=b;
    assign z=c;
    assign y=b;

endmodule
